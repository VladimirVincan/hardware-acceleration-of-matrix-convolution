`ifndef FFT2_DIN_SEQ_LIB_SV
`define FFT2_DIN_SEQ_LIB_SV

`include "din/sequences/fft2_din_base_seq.sv"
`include "din/sequences/fft2_din_simple_seq.sv"
    
`endif