/****************************************************************************
    +-+-+-+-+-+-+-+-+-+-+ +-+-+-+-+-+-+-+-+-+-+-+-+ +-+-+ +-+-+-+-+-+-+-+-+
    |F|u|n|c|t|i|o|n|a|l| |V|e|r|i|f|i|c|a|t|i|o|n| |o|f| |H|a|r|d|w|a|r|e|
    +-+-+-+-+-+-+-+-+-+-+ +-+-+-+-+-+-+-+-+-+-+-+-+ +-+-+ +-+-+-+-+-+-+-+-+

    FILE            fft2_test_lib.sv

    DESCRIPTION     test includes

 ****************************************************************************/

`ifndef FFT2_TEST_LIB_SV
`define FFT2_TEST_LIB_SV

`include "fft2_test_base.sv"
`include "fft2_test_simple.sv"
    
`endif