library verilog;
use verilog.vl_types.all;
entity fft2_pkg is
end fft2_pkg;
