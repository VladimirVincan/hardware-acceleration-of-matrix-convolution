`ifndef CANNY_DIN_SEQ_LIB_SV
`define CANNY_DIN_SEQ_LIB_SV

`include "din/sequences/canny_din_base_seq.sv"
`include "din/sequences/canny_din_simple_seq.sv"
    
`endif