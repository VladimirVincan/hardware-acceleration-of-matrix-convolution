`ifndef CANNY_DOUT_SEQ_LIB_SV
`define CANNY_DOUT_SEQ_LIB_SV

`include "dout/sequences/canny_dout_base_seq.sv"
`include "dout/sequences/canny_dout_simple_seq.sv"
    
`endif