`ifndef FFT2_INIT_SEQ_LIB_SV
`define FFT2_INIT_SEQ_LIB_SV

// `include "init/sequences/fft2_init_base_seq.sv"
// `include "init/sequences/fft2_init_simple_seq.sv"

  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "fft2_init_base_seq.sv"
  `include "fft2_init_simple_seq.sv"

`endif
