library verilog;
use verilog.vl_types.all;
entity fft2_test_top is
end fft2_test_top;
