`ifndef FFT2_DOUT_SEQ_LIB_SV
`define FFT2_DOUT_SEQ_LIB_SV

`include "dout/sequences/fft2_dout_base_seq.sv"
`include "dout/sequences/fft2_dout_simple_seq.sv"
    
`endif